// first timer
module main

fn main() {
	println("Hello World!")
}

// 191224
